module AND_16(out, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16);
	output out;
	input in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16;
	
	assign out = in1 & in2 & in3 & in4 & in5 & in6 & in7 & in8 & in9 & in10 & in11 & in12 & in13 & in14 & in15 & in16;
endmodule 