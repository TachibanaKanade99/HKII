module majority(out, in1, in2);
	output out;
	input in1, in2;
	and (out,in1,in2);
endmodule 